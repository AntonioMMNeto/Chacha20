// SistemaEmbarcadoChaCha20_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcadoChaCha20_tb (
	);

	wire        sistemaembarcadochacha20_inst_clk_bfm_clk_clk;                 // SistemaEmbarcadoChaCha20_inst_clk_bfm:clk -> [SistemaEmbarcadoChaCha20_inst:clk_clk, SistemaEmbarcadoChaCha20_inst_reset_bfm:clk]
	wire  [7:0] sistemaembarcadochacha20_inst_pio_char_in_bfm_conduit_export;  // SistemaEmbarcadoChaCha20_inst_pio_char_in_bfm:sig_export -> SistemaEmbarcadoChaCha20_inst:pio_char_in_export
	wire  [7:0] sistemaembarcadochacha20_inst_pio_char_out_export;             // SistemaEmbarcadoChaCha20_inst:pio_char_out_export -> SistemaEmbarcadoChaCha20_inst_pio_char_out_bfm:sig_export
	wire  [1:0] sistemaembarcadochacha20_inst_pio_ready_in_bfm_conduit_export; // SistemaEmbarcadoChaCha20_inst_pio_ready_in_bfm:sig_export -> SistemaEmbarcadoChaCha20_inst:pio_ready_in_export
	wire  [1:0] sistemaembarcadochacha20_inst_pio_ready_out_export;            // SistemaEmbarcadoChaCha20_inst:pio_ready_out_export -> SistemaEmbarcadoChaCha20_inst_pio_ready_out_bfm:sig_export
	wire        sistemaembarcadochacha20_inst_reset_bfm_reset_reset;           // SistemaEmbarcadoChaCha20_inst_reset_bfm:reset -> SistemaEmbarcadoChaCha20_inst:reset_reset_n

	SistemaEmbarcadoChaCha20 sistemaembarcadochacha20_inst (
		.clk_clk              (sistemaembarcadochacha20_inst_clk_bfm_clk_clk),                 //           clk.clk
		.pio_char_in_export   (sistemaembarcadochacha20_inst_pio_char_in_bfm_conduit_export),  //   pio_char_in.export
		.pio_char_out_export  (sistemaembarcadochacha20_inst_pio_char_out_export),             //  pio_char_out.export
		.pio_ready_in_export  (sistemaembarcadochacha20_inst_pio_ready_in_bfm_conduit_export), //  pio_ready_in.export
		.pio_ready_out_export (sistemaembarcadochacha20_inst_pio_ready_out_export),            // pio_ready_out.export
		.reset_reset_n        (sistemaembarcadochacha20_inst_reset_bfm_reset_reset)            //         reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sistemaembarcadochacha20_inst_clk_bfm (
		.clk (sistemaembarcadochacha20_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm sistemaembarcadochacha20_inst_pio_char_in_bfm (
		.sig_export (sistemaembarcadochacha20_inst_pio_char_in_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 sistemaembarcadochacha20_inst_pio_char_out_bfm (
		.sig_export (sistemaembarcadochacha20_inst_pio_char_out_export)  // conduit.export
	);

	altera_conduit_bfm_0003 sistemaembarcadochacha20_inst_pio_ready_in_bfm (
		.sig_export (sistemaembarcadochacha20_inst_pio_ready_in_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 sistemaembarcadochacha20_inst_pio_ready_out_bfm (
		.sig_export (sistemaembarcadochacha20_inst_pio_ready_out_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sistemaembarcadochacha20_inst_reset_bfm (
		.reset (sistemaembarcadochacha20_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sistemaembarcadochacha20_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
