module chacha(
              input wire           clk,
              input wire           reset_n,
              input wire           read,
              input wire           write,
              input wire [7 : 0]   addr,
              input wire [31 : 0]  write_data,
              output wire [31 : 0] read_data
             );

  //----------------------------------------------------------------
  // Internal constant and parameter definitions.
  //----------------------------------------------------------------
  localparam ADDR_NAME0       = 8'h00;
  localparam ADDR_NAME1       = 8'h01;
  localparam ADDR_VERSION     = 8'h02;

  localparam ADDR_CTRL        = 8'h08;
  localparam CTRL_INIT_BIT    = 0;
  localparam CTRL_NEXT_BIT    = 1;

  localparam ADDR_STATUS      = 8'h09;
  localparam STATUS_READY_BIT = 0;

  localparam ADDR_ROUNDS      = 8'h0b;
  localparam ROUNDS_HIGH_BIT  = 4;
  localparam ROUNDS_LOW_BIT   = 0;

  localparam ADDR_KEY0        = 8'h10;
  localparam ADDR_KEY7        = 8'h17;

  localparam ADDR_IV0         = 8'h20;
  localparam ADDR_IV1         = 8'h21;
  localparam ADDR_IV2         = 8'h22;

  localparam ADDR_DATA_IN0    = 8'h40;
  localparam ADDR_DATA_IN15   = 8'h4f;

  localparam ADDR_DATA_OUT0   = 8'h80;
  localparam ADDR_DATA_OUT15  = 8'h8f;

  localparam CORE_NAME0       = 32'h63686163; // "chac"
  localparam CORE_NAME1       = 32'h68612020; // "ha  "
  localparam CORE_VERSION     = 32'h302e3830; // "0.80"

  localparam DEFAULT_CTR_INIT = 32'h0;


  //----------------------------------------------------------------
  // Registers including update variables and write enable.
  //----------------------------------------------------------------
  reg          init_reg;
  reg          next_reg;
  reg          ctrl_we;

  reg [4 : 0]  rounds_reg;
  reg          rounds_we;

  reg [31 : 0] key_reg [0 : 7];
  reg          key_we;

  reg [31 : 0] iv_reg[0 : 2];
  reg          iv_we;

  reg [31 : 0] data_in_reg [0 : 15];
  reg          data_in_we;


  //----------------------------------------------------------------
  // Wires.
  //----------------------------------------------------------------
  wire [255 : 0] core_key;
  wire [95 : 0]  core_iv;
  wire           core_ready;
  wire [511 : 0] core_data_in;
  wire [511 : 0] core_data_out;
  wire           core_data_out_valid;

  reg [31 : 0]   tmp_read_data;


  //----------------------------------------------------------------
  // Concurrent connectivity for ports etc.
  //----------------------------------------------------------------
  assign core_key     = {key_reg[0], key_reg[1], key_reg[2], key_reg[3],
                         key_reg[4], key_reg[5], key_reg[6], key_reg[7]};

  assign core_iv      = {iv_reg[0], iv_reg[1], iv_reg[2]};

  assign core_data_in = {data_in_reg[00], data_in_reg[01], data_in_reg[02], data_in_reg[03],
                         data_in_reg[04], data_in_reg[05], data_in_reg[06], data_in_reg[07],
                         data_in_reg[08], data_in_reg[09], data_in_reg[10], data_in_reg[11],
                         data_in_reg[12], data_in_reg[13], data_in_reg[14], data_in_reg[15]};

  assign read_data     = tmp_read_data;


  //----------------------------------------------------------------
  // core instantiation.
  //----------------------------------------------------------------
  chacha_core core (
                    .clk(clk),
                    .reset_n(reset_n),
                    .init(init_reg),
                    .next_block(next_reg),
                    .key(core_key),
                    .iv(core_iv),
                    .ctr(DEFAULT_CTR_INIT),
                    .rounds(rounds_reg),
                    .data_in(core_data_in),
                    .ready(core_ready),
                    .data_out(core_data_out),
                    .data_out_valid(core_data_out_valid)
                   );


  //----------------------------------------------------------------
  // reg_update
  //
  // Update functionality for all registers in the core.
  // All registers are positive edge triggered with asynchronous
  // active low reset. All registers have write enable.
  //----------------------------------------------------------------
  always @ (posedge clk)
    begin : reg_update
     integer i;
      if (!reset_n)
        begin
          init_reg   <= 0;
          next_reg   <= 0;
          rounds_reg <= 5'h0;
          iv_reg[0]  <= 32'h0;
          iv_reg[1]  <= 32'h0;
          iv_reg[2]  <= 32'h0;

          for (i = 0 ; i < 8 ; i = i + 1)
            key_reg[i] <= 32'h0;

          for (i = 0 ; i < 16 ; i = i + 1)
            data_in_reg[i] <= 32'h0;
        end
      else
        begin
          if (ctrl_we)
            begin
              init_reg <= write_data[CTRL_INIT_BIT];
              next_reg <= write_data[CTRL_NEXT_BIT];
            end

          if (rounds_we)
            rounds_reg <= write_data[ROUNDS_HIGH_BIT : ROUNDS_LOW_BIT];

          if (key_we)
            key_reg[addr[2 : 0]] <= write_data;

          if (iv_we)
            iv_reg[addr[0]] <= write_data;

          if (data_in_we)
            data_in_reg[addr[3 : 0]] <= write_data;
        end
    end // reg_update


  //----------------------------------------------------------------
  // Address decoder logic.
  //----------------------------------------------------------------
  always @*
    begin : addr_decoder
      ctrl_we       = 0;
      rounds_we     = 0;
      key_we        = 0;
      iv_we         = 0;
      data_in_we    = 0;
      tmp_read_data = 32'h0;


      if (write)
        begin
          if (addr == ADDR_CTRL)
            ctrl_we = 1;

          if (addr == ADDR_ROUNDS)
            rounds_we = 1;

          if ((addr >= ADDR_KEY0) && (addr <= ADDR_KEY7))
            key_we = 1;

          if ((addr >= ADDR_IV0) && (addr <= ADDR_IV2))
            iv_we = 1;

          if ((addr >= ADDR_DATA_IN0) && (addr <= ADDR_DATA_IN15))
            data_in_we = 1;

        end // if (we)

      else if (read)
        begin
          if ((addr >= ADDR_KEY0) && (addr <= ADDR_KEY7))
            tmp_read_data = key_reg[addr[2 : 0]];

          if ((addr >= ADDR_DATA_OUT0) && (addr <= ADDR_DATA_OUT15))
            tmp_read_data = core_data_out[(15 - (addr - ADDR_DATA_OUT0)) * 32 +: 32];

          case (addr)
            ADDR_NAME0:   tmp_read_data = CORE_NAME0;
            ADDR_NAME1:   tmp_read_data = CORE_NAME1;
            ADDR_VERSION: tmp_read_data = CORE_VERSION;
            ADDR_CTRL:    tmp_read_data = {30'h0, next_reg, init_reg};
            ADDR_STATUS:  tmp_read_data = {30'h0, core_data_out_valid, core_ready};
            ADDR_ROUNDS:  tmp_read_data = {27'h0, rounds_reg};
            ADDR_IV0:     tmp_read_data = iv_reg[0];
            ADDR_IV1:     tmp_read_data = iv_reg[1];
            ADDR_IV2:     tmp_read_data = iv_reg[2];

            default:
              begin
              end
          endcase // case (address)
        end
        
    end // addr_decoder
endmodule // chacha
