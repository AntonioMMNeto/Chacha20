
module SistemaEmbarcadoChaChaVerilog (
	clk_clk,
	reset_reset_n);	

	input		clk_clk;
	input		reset_reset_n;
endmodule
